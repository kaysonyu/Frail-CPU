`ifndef __TEST_SVH__
`define __TEST_SVH__


parameter BHT=7;
parameter JHT=4;
parameter RPCT=12;

`endif